module IF_Stage(clk, rst, freeze, Branch_taken, BranchAddr, PC, Instruction);
  input clk, rst, freeze, Branch_taken;
  input[31:0] BranchAddr;
  output[31:0] PC,Instruction;
  
  wire[31:0] InstMemory[63:0];
  wire[31:0] PC_in;
  reg[31:0] PC_out;
  
  always@(posedge clk, posedge rst)
  begin
    if(rst)
      PC_out <= 32'b0;
    else if(freeze) 
      PC_out <= PC_out;
    else
      PC_out <= PC_in;
  end

  assign Instruction = InstMemory[PC_out >>2];
  assign PC = PC_out + 32'd4;
  assign PC_in = (Branch_taken)? BranchAddr: PC;
  
 	assign InstMemory[0] = 32'b11100011101000000000000000010100;
 	assign InstMemory[1] = 32'b11100011101000000001101000000001;
 	assign InstMemory[2] = 32'b11100011101000000010000100000011;
 	assign InstMemory[3] = 32'b11100000100100100011000000000010;
 	assign InstMemory[4] = 32'b11100000101000000100000000000000;
 	assign InstMemory[5] = 32'b11100000010001000101000100000100;
 	assign InstMemory[6] = 32'b11100000110000000110000010100000;
 	assign InstMemory[7] = 32'b11100001100001010111000101000010;
 	assign InstMemory[8] = 32'b11100000000001111000000000000011; 
 	assign InstMemory[9] = 32'b11100001111000001001000000000110;
 	assign InstMemory[10]= 32'b11100000001001001010000000000101;
 	assign InstMemory[11]= 32'b11100001010110000000000000000110; 
 	assign InstMemory[12]= 32'b00010000100000010001000000000001;
 	assign InstMemory[13]= 32'b11100001000110010000000000001000;
 	assign InstMemory[14]= 32'b00000000100000100010000000000010;
 	assign InstMemory[15]= 32'b11100011101000000000101100000001; 
 	assign InstMemory[16]= 32'b11100100100000000001000000000000; 
 	assign InstMemory[17]= 32'b11100100100100001011000000000000;
 	assign InstMemory[18]= 32'b11100100100000000010000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
  assign InstMemory[19]= 32'b11100100100000000011000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
  assign InstMemory[20]= 32'b11100100100000000100000000001100; //STR R4 ,[R0],#13 //MEM[1036] = 41
  assign InstMemory[21]= 32'b11100100100000000101000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
  assign InstMemory[22]= 32'b11100100100000000110000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
  assign InstMemory[23]= 32'b11100100100100001010000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
  assign InstMemory[24]= 32'b11100100100000000111000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
  assign InstMemory[25]= 32'b11100011101000000001000000000100; //MOV R1 ,#4 //R1 = 4
  assign InstMemory[26]= 32'b11100011101000000010000000000000; //MOV R2 ,#0 //R2 = 0
  assign InstMemory[27]= 32'b11100011101000000011000000000000; //MOV R3 ,#0 //R3 = 0
  assign InstMemory[28]= 32'b11100000100000000100000100000011; //ADD R4 ,R0,R3,LSL #2
  assign InstMemory[29]= 32'b11100100100101000101000000000000; //LDR R5 ,[R4],#0
  assign InstMemory[30]= 32'b11100100100101000110000000000100; //LDR R6 ,[R4],#4
  assign InstMemory[31]= 32'b11100001010101010000000000000110; //CMP R5 ,R6
  assign InstMemory[32]= 32'b11000100100001000110000000000000; //STRGT R6 ,[R4],#0
  assign InstMemory[33]= 32'b11000100100001000101000000000100; //STRGT R5 ,[R4],#4
  assign InstMemory[34]= 32'b11100010100000110011000000000001; //ADD R3 ,R3,#1
  assign InstMemory[35]= 32'b11100011010100110000000000000011; //CMP R3 ,#3
  assign InstMemory[36]= 32'b10111010111111111111111111110111; //BLT #-9
  assign InstMemory[37]= 32'b11100010100000100010000000000001; 
  assign InstMemory[38]= 32'b11100001010100100000000000000001; //CMP R2 ,R1
  assign InstMemory[39]= 32'b10111010111111111111111111110011 ; //BLT #-13
  assign InstMemory[40]= 32'b11100100100100000001000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
  assign InstMemory[41]= 32'b11100100100100000010000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
  assign InstMemory[42]= 32'b11100100100100000011000000001000; //STR R3 ,[R0],#8 //R3 = 41
  assign InstMemory[43]= 32'b11100100100100000100000000001100; //STR R4 ,[R0],#12 //R4 = 8192
  assign InstMemory[44]= 32'b11100100100100000101000000010000; //STR R5 ,[R0],#16 //R5 = -123
  assign InstMemory[45]= 32'b11100100100100000110000000010100; //STR R6 ,[R0],#20 //R4 = 10
  assign InstMemory[46]= 32'b11101010111111111111111111111111 ; //B #-1 
 	
endmodule 
      
